// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Thu May 30 20:06:16 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module LEDGcontrol_SM (
    reset,clock,counter[2:0],
    control,counter_reset);

    input reset;
    input clock;
    input [2:0] counter;
    tri0 reset;
    tri0 [2:0] counter;
    output control;
    output counter_reset;
    reg control;
    reg counter_reset;
    reg [1:0] fstate;
    reg [1:0] reg_fstate;
    parameter state1=0,state2=1;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or counter)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            control <= 1'b0;
            counter_reset <= 1'b0;
        end
        else begin
            control <= 1'b0;
            counter_reset <= 1'b0;
            case (fstate)
                state1: begin
                    if ((counter[2:0] == 3'b010))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    control <= 1'b0;

                    if ((counter[2:0] == 3'b100))
                        counter_reset <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        counter_reset <= 1'b0;
                end
                state2: begin
                    if ((counter[2:0] == 3'b100))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    control <= 1'b1;
                end
                default: begin
                    control <= 1'bx;
                    counter_reset <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // LEDGcontrol_SM
